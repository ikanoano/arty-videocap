../vivado-library/ip/dvi2rgb/src/ChannelBond.vhd