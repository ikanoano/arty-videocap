../vivado-library/ip/dvi2rgb/src/SyncBase.vhd