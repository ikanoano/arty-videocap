../ArtyEtherentTX/hdl/ethernet_test.vhd