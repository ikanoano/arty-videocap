../vivado-library/ip/dvi2rgb/src/DVI_Constants.vhd