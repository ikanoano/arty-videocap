../vivado-library/ip/dvi2rgb/src/SyncAsync.vhd