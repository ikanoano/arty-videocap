../vivado-library/ip/dvi2rgb/src/TMDS_Receiver.vhd