../ArtyEtherentTX/hdl/nibble_data.vhd