../ArtyEtherentTX/hdl/add_preamble.vhd