../ArtyEtherentTX/hdl/add_crc32.vhd