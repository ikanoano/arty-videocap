../vivado-library/ip/dvi2rgb/src/InputSERDES.vhd