../vivado-library/ip/dvi2rgb/src/PhaseAlign.vhd